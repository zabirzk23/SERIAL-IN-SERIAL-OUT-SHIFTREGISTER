library verilog;
use verilog.vl_types.all;
entity SISOSR_vlg_vec_tst is
end SISOSR_vlg_vec_tst;
